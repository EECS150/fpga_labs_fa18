module structural_adder (
    input [13:0] a,
    input [13:0] b,
    output [14:0] sum
);
    // Insert your RTL here to create a 14-bit ripple carry adder
    // You will have to use a for-generate loop as outlined in the lab spec
    // Remove this assign statement once you write your own RTL
    assign sum = 15'd0;
endmodule
